module kogg_stone (
	input[15:0] data1, data2,
	output res	
);

endmodule